** sch_path: /home/designer/shared/IPD413_202501/xschem/Tareas/Tarea_1/nmoslv_instrinsic_gain_IPD413-202501-HW1.sch
**.subckt nmoslv_instrinsic_gain_IPD413-202501-HW1 ref g1 d1
*.ipin ref
*.iopin g1
*.iopin d1
E1 g1 GND d1 ref 100
I0 VDD d1 157u
XM1 d1 g1 GND GND sg13_lv_nmos w=120u l=0.5u ng=12 m=1
**** begin user architecture code

*.option wnflag=1
vds ref 0 0.9
vsup VDD 0 1.8

.control
save all

dc vds 0.2 1.8 0.01
plot abs(1/deriv(v(g1)))
*wrdata /home/designer/shared/IPD413_202501_HW1/sim_data/data_nmos_intrinsic_gain_Lp15.dat abs(1/deriv(v(g1)))
wrdata /workspaces/usm-vlsi-tools/shared_xserver/simulations/Projects/IHP/IPD413_2025/sim_data/Tarea_1/data_nmos_intrinsic_gain_Lp15.dat abs(1/deriv(v(g1)))
.endc



.param corner=0

.if (corner==0)
.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ
.endif

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end

** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/simulations/Projects/IHP/IPD413_202501/xschem/Tareas/Tarea_1/nmoslv_charac_IPD413-202501-HW1.sch
**.subckt nmoslv_charac_IPD413-202501-HW1 g1 d1
*.ipin g1
*.iopin d1
XM1 d1 g1 GND GND sg13_lv_nmos w=5u l=0.5u ng=1 m=1
**** begin user architecture code



vgs g1 0 dc=0.75
vds d1 0 dc=0.75

.control
save all
*pre_osdi /home/jmarin/Documents/IHP_designs/ihp_design/psp103_nqs.osdi
*  set color0 = white

save @n.xm1.nsg13_lv_nmos[ids]
save @n.xm1.nsg13_lv_nmos[gm]


*dc vgs 0.01 1.8 0.01
dc vds 0.01 1.8 0.01 vgs 0.1 1.8 0.3

let idn = @n.xm1.nsg13_lv_nmos[ids]
let gmn = @n.xm1.nsg13_lv_nmos[gm]
let vthn = @n.xm1.nsg13_lv_nmos[vth]
let vgsn = @n.xm1.nsg13_lv_nmos[vgs]
let vdsatn = @n.xm1.nsg13_lv_nmos[vdss]
let cgg = @n.xm1.nsg13_lv_nmos[cgg]
let cgsol = @n.xm1.nsg13_lv_nmos[cgsol]
let cgdol = @n.xm1.nsg13_lv_nmos[cgdol]
let vov = 2*idn/gmn
let gmoverId = gmn/idn
let cgg_tot = cgg + cgsol + cgdol
let ft = 1e-9*gmn/6.28/cgg_tot

plot idn
*plot ylog idn
*plot gmn
*plot xlog gmoverId

*wrdata /home/designer/shared/IPD413_202501/sim_data/data_nmos_idvgs_VDSp9_test.txt idn
*wrdata /workspaces/usm-vlsi-tools/shared_xserver/simulations/Projects/IHP/IPD413_202501/sim_data/Tarea_1/data_nmos_idvgs_VDSp9_test.txt idn
wrdata data_nmos_idvgs_VDSp9_test.txt idn

*wrdata /home/designer/shared/IPD413_202501/sim_data/data_nmos_idvgs_VDSp9_gmid-ft.txt gmoverId ft
wrdata data_nmos_idvgs_VDSp9_gmid-ft.txt gmoverId ft

*let W = 5e-6
*setscale gmoverId
*plot idn/W
*plot vov

.endc




.param corner=0

.if (corner==0)
.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ
.endif

**** end user architecture code
**.ends
.GLOBAL GND
.end

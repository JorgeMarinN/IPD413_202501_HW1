** sch_path: /home/designer/shared/IPD413_202501_HW1/nmoslv_charac_IPD413-202501-HW1.sch
**.subckt nmoslv_charac_IPD413-202501-HW1 g1 d1
*.ipin g1
*.iopin d1
XM1 d1 g1 GND GND sg13_lv_nmos w=5u l=0.5u ng=1 m=1
**** begin user architecture code



vgs g1 0 dc=0.9
vds d1 0 dc=0.9

.control
save all
*pre_osdi /home/jmarin/Documents/IHP_designs/ihp_design/psp103_nqs.osdi
*  set color0 = white

save @n.xm1.nsg13_lv_nmos[ids]
save @n.xm1.nsg13_lv_nmos[gm]


dc vgs 0.01 1.8 0.01

let idn = @n.xm1.nsg13_lv_nmos[ids]
let gmn = @n.xm1.nsg13_lv_nmos[gm]
let vthn = @n.xm1.nsg13_lv_nmos[vth]
let vgsn = @n.xm1.nsg13_lv_nmos[vgs]
let vdsatn = @n.xm1.nsg13_lv_nmos[vdss]
let vov1 = v(g1) - vthn
let vov2 = 2*idn/gmn
let gmoverId = gmn/idn

plot idn
*plot idn vs vov1
*plot idn vs vov2
*plot vov2
plot gmn
plot xlog gmoverId
*plot idn vs vdsatn

let W = 5e-6
*let gmoverId = gmn/idn
setscale gmoverId
plot idn/W
plot vov2



*wrdata /foss/designs/UNIC-CASS_OS_analog_flow/data_nmos_idvgs_VDSp9_test.txt idn


.endc




.param corner=0

.if (corner==0)
.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ
.endif

**** end user architecture code
**.ends
.GLOBAL GND
.end

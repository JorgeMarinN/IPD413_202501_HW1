** sch_path: /home/designer/shared/IPD413_202501/xschem/Tareas/Tarea_1/cs_amp_full_IPD413HW1.sch
**.subckt cs_amp_full_IPD413HW1 ref g1 d1 g2 vout
*.ipin ref
*.iopin g1
*.iopin d1
*.iopin g2
*.iopin vout
E1 g1 GND d1 ref 1000
I0 VDD d1 157u
I1 VDD vout 157u
XM1 d1 g1 GND GND sg13_lv_nmos w=120u l=0.5u ng=12 m=1
XM2 vout g2 GND GND sg13_lv_nmos w=120u l=0.5u ng=12 m=1
**** begin user architecture code

.option wnflag=1
vds ref 0 0.9
vsup VDD 0 1.8
vin g1 g2 dc=0 ac=1

cload vout 0 5p

.control
save all

save @m.xm2.msky130_fd_pr__nfet_01v8[gm]
save @m.xm2.msky130_fd_pr__nfet_01v8[id]
save @m.xm2.msky130_fd_pr__nfet_01v8[gds]

dc vin -0.01 0.01 0.001

let gdsn = @m.xm2.msky130_fd_pr__nfet_01v8[gds]
let gmn = @m.xm2.msky130_fd_pr__nfet_01v8[gm]
let idn = @m.xm2.msky130_fd_pr__nfet_01v8[id]
let ao = gmn / gdsn

plot deriv(v(vout)) vs v(vout) ao vs v(vout)

ac dec 100 1 1T
plot vdb(vout)

.endc



.param corner=0

.if (corner==0)
.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ
.endif

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
